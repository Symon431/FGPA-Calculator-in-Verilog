library verilog;
use verilog.vl_types.all;
entity tb_adder_subtractor is
end tb_adder_subtractor;
