module adder_subtractor (
    input [3:0] A,
    input [3:0] B,
    input OP,  // 0 = add, 1 = subtract
    output [7:0] S
);

    wire [3:0] B_muxed;
    wire [3:0] Sum;
    wire Cout;
    wire Cin;

    // Choose between B and ~B. So if OP value is 0 B_muxed will be B and if its 1(subtraction) it will be ~B 
    mux2to1 B_selector (
        .in0(B),
        .in1(~B),
        .sel(OP),
        .out(B_muxed)
    );

    // Choose Cin = 0 (add) or 1 (sub)
    mux2to1_1bit Cin_selector (
        .in0(1'b0),
        .in1(1'b1),
        .sel(OP),
        .out(Cin)
    );

    // Perform the actual addition/subtraction
    ripple_carry_adder_4bit RCA (
        .A(A),
        .B(B_muxed),
        .Cin(Cin),
        .Sum(Sum),
        .Cout(Cout)
    );

    // Output: pad 3 zeros, then Cout and Sum
    assign S = {3'b000, Cout, Sum};

endmodule

