module ripple_carry_adder_4bit (
    input [3:0] A,
    input [3:0] B,
    input Cin,
    output [3:0] Sum,
    output Cout
);

    wire c1, c2, c3; // internal carry wires

    // Instantiate four 1-bit full adders
    full_adder_1bit fa0 (
        .A(A[0]),
        .B(B[0]),
        .Cin(Cin),
        .Sum(Sum[0]),
        .Cout(c1)
    );

    full_adder_1bit fa1 (
        .A(A[1]),
        .B(B[1]),
        .Cin(c1),
        .Sum(Sum[1]),
        .Cout(c2)
    );

    full_adder_1bit fa2 (
        .A(A[2]),
        .B(B[2]),
        .Cin(c2),
        .Sum(Sum[2]),
        .Cout(c3)
    );

    full_adder_1bit fa3 (
        .A(A[3]),
        .B(B[3]),
        .Cin(c3),
        .Sum(Sum[3]),
        .Cout(Cout)
    );

endmodule



module mux2to1_1bit (
    input in0,
    input in1,
    input sel,
    output out
);
    assign out = sel ? in1 : in0;
endmodule



module mux2to1 (
    input [3:0] in0,
    input [3:0] in1,
    input sel,
    output [3:0] out
);
    assign out = sel ? in1 : in0;
endmodule



module full_adder_1bit (
    input A, B, Cin,
    output reg Sum, Cout
);

always @(*) begin
    {Cout, Sum} = A + B + Cin;  
end

endmodule


module fsm (
    input clk,
    input reset,
    input start,
    input enter,

    output reg [2:0] op_code,      // Controls datapath (LOAD_A, COMPUTE, etc.)
    output reg wrt_addr,           // Selects register A or B
    output reg [1:0] compute_op,   // Operation selection (passed from top level)
    output reg [2:0] state         // Current FSM state (for HEX3 display)
);

    // FSM State Encoding
    localparam IDLE     = 3'b000,
               START    = 3'b001,
               GET_A    = 3'b010,
               DISP_A   = 3'b011,
               GET_B    = 3'b100,
               DISP_B   = 3'b101,
               COMPUTE  = 3'b110,
               RESULT   = 3'b111;

    reg [2:0] next_state;

    // Sequential logic: state transition
    always @(posedge clk or posedge reset) begin
        if (reset)
            state <= IDLE;
        else
            state <= next_state;
    end

    // Combinational logic: next state + control outputs
    always @(*) begin
        // Default values
        op_code = 3'b000;       // NOOP
        wrt_addr = 0;
        compute_op = 2'b00;
        next_state = state;

        case (state)
            IDLE: begin
                if (start)
                    next_state = START;
            end

            START: begin
                op_code = 3'b111;       // RESET (optional)
                next_state = GET_A;
            end

            GET_A: begin
                wrt_addr = 0;           // Select reg_A
                if (enter)
                    next_state = DISP_A;
            end

            DISP_A: begin
                op_code = 3'b010;       // DISPLAY_A
                if (!enter)
                    next_state = GET_B;
            end

            GET_B: begin
                wrt_addr = 1;           // Select reg_B
                if (enter)
                    next_state = DISP_B;
            end

            DISP_B: begin
                op_code = 3'b100;       // DISPLAY_B
                if (!enter)
                    next_state = COMPUTE;
            end

            COMPUTE: begin
                op_code = 3'b101;       // COMPUTE
                // `compute_op` will be driven by top-level and passed through in datapath
                next_state = (enter) ? RESULT : COMPUTE;
            end

            RESULT: begin
                op_code = 3'b110;       // DISPLAY_RESULT
                next_state = IDLE;
            end
        endcase
    end

endmodule





module display_logic (
    input  wire [7:0] binary_in,
    output reg  [6:0] seg_hundreds,
    output reg  [6:0] seg_tens,
    output reg  [6:0] seg_ones
);

    reg [3:0] hundreds, tens, ones;

    always @(*) begin
        hundreds = binary_in / 100;
        tens     = (binary_in % 100) / 10;
        ones     = binary_in % 10;

        // Hundreds
        case (hundreds)
            4'd0: seg_hundreds = 7'b1000000;
            4'd1: seg_hundreds = 7'b1111001;
            4'd2: seg_hundreds = 7'b0100100;
            4'd3: seg_hundreds = 7'b0110000;
            4'd4: seg_hundreds = 7'b0011001;
            4'd5: seg_hundreds = 7'b0010010;
            4'd6: seg_hundreds = 7'b0000010;
            4'd7: seg_hundreds = 7'b1111000;
            4'd8: seg_hundreds = 7'b0000000;
            4'd9: seg_hundreds = 7'b0010000;
            default: seg_hundreds = 7'b1111111;
        endcase

        // Tens
        case (tens)
            4'd0: seg_tens = 7'b1000000;
            4'd1: seg_tens = 7'b1111001;
            4'd2: seg_tens = 7'b0100100;
            4'd3: seg_tens = 7'b0110000;
            4'd4: seg_tens = 7'b0011001;
            4'd5: seg_tens = 7'b0010010;
            4'd6: seg_tens = 7'b0000010;
            4'd7: seg_tens = 7'b1111000;
            4'd8: seg_tens = 7'b0000000;
            4'd9: seg_tens = 7'b0010000;
            default: seg_tens = 7'b1111111;
        endcase

        // Ones
        case (ones)
            4'd0: seg_ones = 7'b1000000;
            4'd1: seg_ones = 7'b1111001;
            4'd2: seg_ones = 7'b0100100;
            4'd3: seg_ones = 7'b0110000;
            4'd4: seg_ones = 7'b0011001;
            4'd5: seg_ones = 7'b0010010;
            4'd6: seg_ones = 7'b0000010;
            4'd7: seg_ones = 7'b1111000;
            4'd8: seg_ones = 7'b0000000;
            4'd9: seg_ones = 7'b0010000;
            default: seg_ones = 7'b1111111;
        endcase
    end

endmodule



module calculator_datapath (
    input clk,
    input reset,
    input [3:0] data_in,
    input [2:0] op_code,         // Instruction: LOAD A, LOAD B, COMPUTE, etc.
    input [1:0] compute_op,      // Operation for ALU: ADD, SUB, etc.
    output [7:0] result,
    output done,
    output negative,
    output div_by_zero
);

    // Derived control signals
    wire load_signal = (op_code == 3'b001 || op_code == 3'b011); // LOAD A or B
    wire write_addr  = op_code[1];  // 0 for A (001), 1 for B (011)
    wire [1:0] sel;                 // Load signals to reg_A and reg_B

    // Register outputs
    wire [3:0] A, B;

    // Decoder to select which register to load
    decoder_1to2 dec (
        .write_addr(write_addr),
        .load(load_signal),
        .sel(sel)
    );

    // Register A (load when sel[0] is 1)
    dff4 reg_A (
        .clk(clk),
        .reset(reset),
        .load(sel[0]),
        .d(data_in),
        .q(A)
    );

    // Register B (load when sel[1] is 1)
    dff4 reg_B (
        .clk(clk),
        .reset(reset),
        .load(sel[1]),
        .d(data_in),
        .q(B)
    );

    // ALU (computes and outputs final result)
    alu alu_inst (
        .clk(clk),
        .reset(reset),
        .A(A),
        .B(B),
        .op_code(op_code),
        .compute_op(compute_op),
        .result(result),
        .done(done),
        .div_by_zero(div_by_zero),
        .negative(negative)
    );

endmodule



module calculator (
    input clk,
    input reset,
    input start,
    input enter,
    input [3:0] data_in,
    input [2:0] op_code,
    input [1:0] compute_op,
    output [6:0] HEX0, HEX1, HEX2,
    output [2:0] HEX3,
    output [7:0] result,           
    output done, negative, div_by_zero
);

    wire [2:0] state;
    wire [7:0] result_internal;

    // FSM to control instruction entry flow
    fsm fsm_inst (
        .clk(clk),
        .reset(reset),
        .start(start),
        .enter(enter),
        .state(state)
    );

    // Datapath to execute instructions
    calculator_datapath dp (
        .clk(clk),
        .reset(reset),
        .data_in(data_in),
        .op_code(op_code),
        .compute_op(compute_op),
        .result(result_internal),     // internal wire
        .done(done),
        .negative(negative),
        .div_by_zero(div_by_zero)
    );

    // Display logic for converting binary to BCD segments
    display_logic display (
        .binary_in(result_internal),
        .seg_hundreds(HEX2),
        .seg_tens(HEX1),
        .seg_ones(HEX0)
    );

    assign HEX3 = state;
    assign result = result_internal;  

endmodule


module dff4 (
    input clk,
    input reset,
    input load,             // Enables writing into register
    input [3:0] d,          // Input data
    output reg [3:0] q      // Stored output
);

    always @(posedge clk or posedge reset) begin
        if (reset)
            q <= 4'b0000;
        else if (load)
            q <= d;
    end

endmodule

//The calculator needs two 4-bit registers (reg_A and reg_B) to hold input numbers before computation. The module comes into play



module decoder_1to2 (
    input write_addr,       // 0 ? A, 1 ? B
    input load,             // Enable loading
    output reg [1:0] sel    //The output(select line) - depends on the value of write_adder(selector)
);

    always @(*) begin
        if (load) begin
            sel = (write_addr == 1'b0) ? 2'b01 : 2'b10;  
        end else begin
            sel = 2'b00;
        end
    end

endmodule




module alu (
    input clk,
    input reset,
    input [3:0] A,
    input [3:0] B,
    input [2:0] op_code,       // Main instruction code
    input [1:0] compute_op,    // Specific compute operation: ADD, SUB, MUL, DIV
    output reg [7:0] result,   // 8-bit result
    output reg done,           // Operation complete flag
    output reg div_by_zero,    // Division-by-zero flag
    output reg negative        // Negative result flag (subtraction only)
);

    // Intermediate result from adder-subtractor
    wire [7:0] add_sub_result;

    // Adder-Subtractor instance (matches current definition)
    adder_subtractor add_sub (
        .A(A),
        .B(B),
        .OP(compute_op[0]),  // 0 = ADD, 1 = SUB
        .S(add_sub_result)   // Result is {3'b000, Cout, Sum}
    );

    always @(posedge clk or posedge reset) begin
        if (reset) begin
            result <= 8'b0;
            done <= 0;
            div_by_zero <= 0;
            negative <= 0;
        end else begin
            done <= 0;
            div_by_zero <= 0;
            negative <= 0;

            case (op_code)
                3'b101: begin // COMPUTE
                    case (compute_op)
                        2'b00: begin
                            result <= add_sub_result; // ADD
                            done <= 1;
                        end
                      
                      2'b01: begin
                        done <= 1;
                          if (A >= B)
                            result <= {4'b0000, A - B};
                          else begin
                            result <= {4'b0000, B - A};
                            negative <= 1;
                        end
                      end

                        2'b11: begin
                            if (B == 0) begin
                                div_by_zero <= 1;
                                result <= 8'b0;
                            end else begin
                                result <= {A % B, A / B};
                                done <= 1;
                            end
                        end
                        
                        
                        2'b10: begin
                       // MUL
                        result <= A * B;
                          done <= 1;
                      end
                        
                        
                    endcase
                end
                
                      

                3'b010: begin // DISPLAY A
                    result <= {4'b0000, A};
                    done <= 1;
                end

                3'b100: begin // DISPLAY B
                    result <= {4'b0000, B};
                    done <= 1;
                end

                3'b110: begin // DISPLAY RESULT (no update)
                    done <= 1;
                end

                3'b000: begin // NOOP
                    done <= 0;
                end

                default: begin
                    done <= 0;
                    div_by_zero <= 0;
                    negative <= 0;
                end
            endcase
        end
    end
endmodule




module adder_subtractor (
    input [3:0] A,
    input [3:0] B,
    input OP,  // 0 = add, 1 = subtract
    output [7:0] S
);

    wire [3:0] B_muxed;
    wire [3:0] Sum;
    wire Cout;
    wire Cin;

    // Choose between B and ~B. So if OP value is 0 B_muxed will be B and if its 1(subtraction) it will be ~B 
    mux2to1 B_selector (
        .in0(B),
        .in1(~B),
        .sel(OP),
        .out(B_muxed)
    );

    // Choose Cin = 0 (add) or 1 (sub)
    mux2to1_1bit Cin_selector (
        .in0(1'b0),
        .in1(1'b1),
        .sel(OP),
        .out(Cin)
    );

    // Perform the actual addition/subtraction
    ripple_carry_adder_4bit RCA (
        .A(A),
        .B(B_muxed),
        .Cin(Cin),
        .Sum(Sum),
        .Cout(Cout)
    );

    // Output: pad 3 zeros, then Cout and Sum
    assign S = {4'b0000, Sum};

endmodule






