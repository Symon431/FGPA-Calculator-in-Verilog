library verilog;
use verilog.vl_types.all;
entity tb_dff4 is
end tb_dff4;
