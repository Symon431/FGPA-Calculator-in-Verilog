library verilog;
use verilog.vl_types.all;
entity adder_subtractor is
    port(
        A               : in     vl_logic_vector(3 downto 0);
        B               : in     vl_logic_vector(3 downto 0);
        OP              : in     vl_logic;
        S               : out    vl_logic_vector(7 downto 0)
    );
end adder_subtractor;
