library verilog;
use verilog.vl_types.all;
entity binary_multiplierTB is
end binary_multiplierTB;
