library verilog;
use verilog.vl_types.all;
entity tb_mux2to1 is
end tb_mux2to1;
