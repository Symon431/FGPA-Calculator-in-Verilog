library verilog;
use verilog.vl_types.all;
entity project1b_tb is
end project1b_tb;
