library verilog;
use verilog.vl_types.all;
entity tb_calculator_datapath is
end tb_calculator_datapath;
