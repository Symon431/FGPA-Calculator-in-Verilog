library verilog;
use verilog.vl_types.all;
entity tb_decoder_1to2 is
end tb_decoder_1to2;
