library verilog;
use verilog.vl_types.all;
entity tb_ripple_carry_adder is
end tb_ripple_carry_adder;
